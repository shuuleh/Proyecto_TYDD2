library verilog;
use verilog.vl_types.all;
entity Control1_vlg_vec_tst is
end Control1_vlg_vec_tst;
