-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 06 15:55:28 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Control IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SI_SD : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        D_I : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        PD_PI : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END Control;

ARCHITECTURE BEHAVIOR OF Control IS
    TYPE type_fstate IS (R,D,I,A);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= R;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,SI_SD)
    BEGIN
        D_I <= "0000";
        PD_PI <= "0000";
        CASE fstate IS
            WHEN R =>
                IF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= D;
                ELSIF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= A;
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= I;
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= R;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= R;
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    PD_PI <= "1111";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    PD_PI <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    PD_PI <= "0000";
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    D_I <= "1010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    D_I <= "0010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    D_I <= "1000";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    D_I <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    D_I <= "0000";
                END IF;
            WHEN D =>
                IF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= I;
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= R;
                ELSIF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= A;
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= D;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= D;
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    PD_PI <= "1111";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    PD_PI <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    PD_PI <= "0000";
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    D_I <= "1010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    D_I <= "0010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    D_I <= "1000";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    D_I <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    D_I <= "0000";
                END IF;
            WHEN I =>
                IF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= D;
                ELSIF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= A;
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= R;
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= I;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= I;
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    PD_PI <= "1111";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    PD_PI <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    PD_PI <= "0000";
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    D_I <= "1010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    D_I <= "0010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    D_I <= "1000";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    D_I <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    D_I <= "0000";
                END IF;
            WHEN A =>
                IF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= I;
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= R;
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= D;
                ELSIF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= A;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= A;
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    PD_PI <= "1111";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    PD_PI <= "0101";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    PD_PI <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    PD_PI <= "0000";
                END IF;

                IF ((SI_SD(1 DOWNTO 0) = "00")) THEN
                    D_I <= "1010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "01")) THEN
                    D_I <= "0010";
                ELSIF ((SI_SD(1 DOWNTO 0) = "10")) THEN
                    D_I <= "1000";
                ELSIF ((SI_SD(1 DOWNTO 0) = "11")) THEN
                    D_I <= "0101";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    D_I <= "0000";
                END IF;
            WHEN OTHERS => 
                D_I <= "XXXX";
                PD_PI <= "XXXX";
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
