library verilog;
use verilog.vl_types.all;
entity TyDD_vlg_vec_tst is
end TyDD_vlg_vec_tst;
